
module ifu(
    input clk_i,
    output [31:0] pc_o,
    input [31:0] instr_in,
    output [31:0] instr_out
);

    reg [31:0] pc_r;
    


endmodule