module pipe_exu import liang_pkg::*;
(
  input logic clk_i,
  input logic rst_i,
  input logic id_valid_i,
  input idToEx_t idToEx_i,
  output logic ex_ready_o,

  output logic ex_valid_o,
  output exToWb_t exToWb_o 
);

  



endmodule