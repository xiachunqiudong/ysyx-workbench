module inst_buffer
(
  input clk_i,
  input rst_i
);




endmodule
