module fifo(
  input logic1 clk,
  input data_in,
  output data_out,
  output logic empty_o,
  output logic full_o
);

endmodule