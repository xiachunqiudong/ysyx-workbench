module ifu_icache_data_array(
  input clk_i
);

endmodule